/*******************************************************************
 *
 * ETF Comment header
 *
 *******************************************************************/
/*******************************************************************
 *
 * F = ~D & (A | B | C)
 *
 *******************************************************************/

/*******************************************************************/
module or_3_gate(input i_A, input i_B, input i_C, output o_Y);
    assign o_Y = i_A | i_B | i_C;
endmodule : or_3_gate
/*******************************************************************/

/*******************************************************************/
module inv(input i_A, output o_Y);
    assign o_Y = ~i_A;
endmodule : inv
/*******************************************************************/

/*******************************************************************/
module and_2_gate(input i_A, input i_B, output o_Y);
    assign o_Y = i_A & i_B;
endmodule : and_2_gate
/*******************************************************************/

/*******************************************************************/
module example_1_gate(
    input i_A,
    input i_B,
    input i_C,
    input i_D,
    output [7 : 0] o_Y
);
    
    wire w_x1;
    wire w_not_d;
    wire w_y;
    
    or_3_gate or_3_gate_inst(.i_A(i_A), .i_B(i_B), .i_C(i_C), .o_Y(w_x1));
    
    inv inv_inst(.i_A(i_D), .o_Y(w_not_d));
    
    and_2_gate and_2_gate_inst(.i_A(w_x1), .i_B(w_not_d), .o_Y(w_y));
    
    assign o_Y = {7'h0, w_y};

endmodule : example_1_gate
/*******************************************************************/

