/*******************************************************************
 *
 * ETF Comment header
 *
 *******************************************************************/

/*******************************************************************
 *
 * Logic gate: AND -> Y = A & B
 *  
 *     -------------
 *     | A | B | Y |
 *     -------------
 *     | 0 | 0 | 0 |
 *     -------------
 *     | 0 | 1 | 0 |
 *     -------------
 *     | 1 | 0 | 0 |
 *     -------------
 *     | 1 | 1 | 1 |
 *     -------------
 *
 *******************************************************************/
module and_gate(
    input i_A, 
    input i_B, 
    output o_Y
);
    /** \TODO: Ovdje unijeti logicku funkciju!!! */
	assign o_Y = i_A & i_B;
    
endmodule

